magic
tech scmos
timestamp 1606577988
<< nwell >>
rect -15 2 44 20
<< polysilicon >>
rect -6 8 -4 11
rect 16 8 18 11
rect 36 8 38 11
rect -6 -3 -4 4
rect 16 -1 18 4
rect 36 -1 38 4
rect -5 -9 -4 -3
rect 17 -7 18 -1
rect 37 -7 38 -1
rect -6 -20 -4 -9
rect 16 -20 18 -7
rect 36 -20 38 -7
rect -6 -30 -4 -26
rect 16 -30 18 -26
rect 36 -30 38 -26
<< ndiffusion >>
rect -15 -21 -6 -20
rect -10 -26 -6 -21
rect -4 -26 0 -20
rect 5 -26 16 -20
rect 18 -26 23 -20
rect 29 -26 36 -20
rect 38 -26 39 -20
<< pdiffusion >>
rect -9 4 -6 8
rect -4 4 16 8
rect 18 4 36 8
rect 38 4 40 8
<< metal1 >>
rect -8 14 4 19
rect -13 8 -9 14
rect -13 -9 -10 -3
rect 9 -7 12 -1
rect 30 -7 33 -1
rect 40 -13 44 4
rect 0 -17 44 -13
rect 0 -20 5 -17
rect 39 -20 44 -17
rect -15 -32 -10 -26
rect 23 -32 29 -26
rect -10 -38 -3 -32
rect 3 -38 23 -32
rect 29 -38 40 -32
<< ntransistor >>
rect -6 -26 -4 -20
rect 16 -26 18 -20
rect 36 -26 38 -20
<< ptransistor >>
rect -6 4 -4 8
rect 16 4 18 8
rect 36 4 38 8
<< polycontact >>
rect -10 -9 -5 -3
rect 12 -7 17 -1
rect 33 -7 37 -1
<< ndcontact >>
rect -15 -26 -10 -21
rect 0 -26 5 -20
rect 23 -26 29 -20
rect 39 -26 44 -20
<< pdcontact >>
rect -13 4 -9 8
rect 40 4 44 8
<< psubstratepcontact >>
rect -15 -38 -10 -32
rect -3 -38 3 -32
rect 23 -38 29 -32
<< nsubstratencontact >>
rect -13 14 -8 19
rect 4 14 9 19
<< labels >>
rlabel metal1 -12 -7 -12 -7 3 a
rlabel metal1 10 -4 10 -4 1 b
rlabel metal1 31 -4 31 -4 1 c
rlabel metal1 42 -15 42 -15 7 f
rlabel metal1 -7 -35 -7 -35 1 Gnd
rlabel metal1 -6 16 -6 16 5 Vdd
<< end >>
