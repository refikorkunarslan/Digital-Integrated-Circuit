* SPICE3 file created from nor2.ext - technology: scmos

M1000 a_n4_4# a Vdd Vdd pmos w=4u l=2u
+  ad=80p pd=48u as=28p ps=22u
M1001 f b a_n4_4# Vdd pmos w=4u l=2u
+  ad=60p pd=38u as=0p ps=0u
M1002 f a Gnd Gnd nmos w=6u l=2u
+  ad=120p pd=52u as=186p ps=86u
M1003 Gnd b f Gnd nmos w=6u l=2u
+  ad=0p pd=0u as=0p ps=0u
C0 Vdd a 1.7fF
C1 Vdd b 1.7fF
C2 Vdd f 0.5fF
C3 b f 0.3fF
C4 Gnd Gnd 13.5fF
C5 f Gnd 10.1fF
C6 b  Gnd 9.1fF
C7 a Gnd  9.1fF

VCC    Vdd     Gnd     DC=2.5


* The following two lines are for TRANSIENT analysis
*
*Vname +Node -Node Option T1  V1   T2  V2   T3   V3    T4  V4  T5   V5 
*----- ----- ----- ------ --  --   --  --   ---- --    --  --  ---- -- 
Vin     a     f    PWL(   0   0    4N  0    4.1N 2.5   8N  2.5 8.1N  0  ) 

* The following two lines are for TRANSIENT analysis
*
*Vname +Node -Node Option T1  V1   T2  V2   T3   V3    T4  V4  T5   V5 
*----- ----- ----- ------ --  --   --  --   ---- --    --  --  ---- -- 
Vi     b     f    PWL(   0   0    4N  0    4.1N 2.5   8N  2.5 8.1N  0  ) 

*     TSTEP TSTOP
*     ----- -----
.TRAN 0.1N  12N


* The following line is for DC analysis

.DC VIN 0 2.6 0.1


* TEMPERATURE and OPTIONS SETTING

.OPTIONS TEMP=25 reltol = 1e-6 

*MODELS

.include tsmc_cmos025

.END
