magic
tech scmos
timestamp 1606574185
<< nwell >>
rect -15 2 34 20
<< polysilicon >>
rect -6 8 -4 11
rect 16 8 18 11
rect -6 -3 -4 4
rect 16 -1 18 4
rect -5 -9 -4 -3
rect 17 -7 18 -1
rect -6 -20 -4 -9
rect 16 -20 18 -7
rect -6 -30 -4 -26
rect 16 -30 18 -26
<< ndiffusion >>
rect -15 -21 -6 -20
rect -10 -26 -6 -21
rect -4 -24 1 -20
rect 6 -24 16 -20
rect -4 -26 16 -24
rect 18 -25 32 -20
rect 38 -25 40 -20
rect 18 -26 40 -25
<< pdiffusion >>
rect -9 4 -6 8
rect -4 4 16 8
rect 18 4 22 8
rect 27 4 33 8
<< metal1 >>
rect -9 15 0 20
rect 5 15 32 20
rect -13 8 -9 15
rect -13 -9 -10 -3
rect 9 -7 12 -1
rect 22 -13 27 4
rect 1 -18 29 -13
rect 1 -20 6 -18
rect -15 -32 -10 -26
rect 32 -32 38 -25
rect -15 -38 -3 -32
rect 3 -38 8 -32
rect 14 -38 32 -32
rect 38 -38 40 -32
<< ntransistor >>
rect -6 -26 -4 -20
rect 16 -26 18 -20
<< ptransistor >>
rect -6 4 -4 8
rect 16 4 18 8
<< polycontact >>
rect -10 -9 -5 -3
rect 12 -7 17 -1
<< ndcontact >>
rect -15 -26 -10 -21
rect 1 -24 6 -20
rect 32 -25 38 -20
<< pdcontact >>
rect -13 4 -9 8
rect 22 4 27 8
<< psubstratepcontact >>
rect -3 -38 3 -32
rect 8 -38 14 -32
rect 32 -38 38 -32
<< nsubstratencontact >>
rect -13 15 -9 20
rect 0 15 5 20
<< labels >>
rlabel metal1 -12 -7 -12 -7 3 a
rlabel metal1 10 -4 10 -4 1 b
rlabel metal1 -9 -36 -9 -36 1 Gnd
rlabel metal1 28 -16 28 -16 1 f
rlabel metal1 -6 17 -6 17 5 Vdd
<< end >>
