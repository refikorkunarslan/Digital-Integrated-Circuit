* SPICE3 file created from nand3.ext - technology: scmos

M1000 f a Vdd Vdd pmos w=4u l=2u
+  ad=104p pd=68u as=104p ps=68u
M1001 Vdd b f Vdd pmos w=4u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1002 f c Vdd Vdd pmos w=4u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1003 a_n4_n26# a Gnd Gnd nmos w=6u l=2u
+  ad=120p pd=52u as=54p ps=30u
M1004 a_18_n26# b a_n4_n26# Gnd nmos w=6u l=2u
+  ad=108p pd=48u as=0p ps=0u
M1005 f c a_18_n26# Gnd nmos w=6u l=2u
+  ad=36p pd=24u as=0p ps=0u
C0 c f 0.3fF
C1 b f 0.3fF
C2 Vdd c 1.7fF
C3 Vdd f 0.8fF
C4 Vdd b 1.7fF
C5 Vdd a 1.7fF
C6 Gnd Gnd 11.8fF
C7 f Gnd 16.0fF
C8 c Gnd 8.7fF
C9 b Gnd 9.1fF
C10 a Gnd 9.1fF

VCC    Vdd     Gnd     DC=2.5


* The following two lines are for TRANSIENT analysis
*
*Vname +Node -Node Option T1  V1   T2  V2   T3   V3    T4  V4  T5   V5 
*----- ----- ----- ------ --  --   --  --   ---- --    --  --  ---- -- 
Vin     a     f    PWL(   0   0    4N  0    4.1N 2.5   8N  2.5 8.1N  0  ) 

* The following two lines are for TRANSIENT analysis
*
*Vname +Node -Node Option T1  V1   T2  V2   T3   V3    T4  V4  T5   V5 
*----- ----- ----- ------ --  --   --  --   ---- --    --  --  ---- -- 
Vi     b     f    PWL(   0   0    4N  0    4.1N 2.5   8N  2.5 8.1N  0  ) 

* The following two lines are for TRANSIENT analysis
*
*Vname +Node -Node Option T1  V1   T2  V2   T3   V3    T4  V4  T5   V5 
*----- ----- ----- ------ --  --   --  --   ---- --    --  --  ---- -- 
V     c     f    PWL(   0   0    4N  0    4.1N 2.5   8N  2.5 8.1N  0  ) 

*     TSTEP TSTOP
*     ----- -----
.TRAN 0.1N  12N


* The following line is for DC analysis

.DC VIN 0 2.6 0.1


* TEMPERATURE and OPTIONS SETTING

.OPTIONS TEMP=25 reltol = 1e-6 

*MODELS

.include tsmc_cmos025

.END
