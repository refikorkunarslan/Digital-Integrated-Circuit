magic
tech scmos
timestamp 1611333839
<< nwell >>
rect 1245 1821 1300 1853
rect 1355 1844 1430 1848
rect 1185 1799 1223 1820
rect 1354 1818 1430 1844
rect 1448 1830 1505 1854
rect 1247 1731 1303 1755
rect 1380 1686 1446 1713
rect 866 1478 922 1502
rect 1239 1489 1294 1521
rect 1349 1512 1432 1516
rect 1348 1490 1432 1512
rect 1765 1494 1821 1518
rect 1179 1467 1217 1488
rect 1348 1486 1431 1490
rect 1031 1417 1127 1441
rect 1241 1399 1297 1423
rect 871 1355 927 1379
rect 1374 1354 1440 1381
rect 867 1199 963 1223
<< ntransistor >>
rect 1260 1797 1262 1803
rect 1282 1797 1284 1803
rect 1468 1820 1470 1823
rect 1199 1789 1201 1792
rect 1374 1794 1376 1800
rect 1396 1794 1398 1800
rect 1261 1705 1263 1711
rect 1283 1705 1285 1711
rect 1400 1662 1402 1668
rect 1422 1662 1424 1668
rect 1254 1465 1256 1471
rect 1276 1465 1278 1471
rect 1779 1468 1781 1474
rect 1801 1468 1803 1474
rect 1849 1468 1851 1473
rect 880 1452 882 1458
rect 902 1452 904 1458
rect 1193 1457 1195 1460
rect 1368 1462 1370 1468
rect 1390 1462 1392 1468
rect 1045 1391 1047 1397
rect 1067 1391 1069 1397
rect 1093 1391 1096 1397
rect 1255 1373 1257 1379
rect 1277 1373 1279 1379
rect 885 1329 887 1335
rect 907 1329 909 1335
rect 1394 1330 1396 1336
rect 1416 1330 1418 1336
rect 825 1173 827 1178
rect 881 1173 883 1179
rect 903 1173 905 1179
rect 929 1173 932 1179
rect 1370 1109 1373 1118
<< ptransistor >>
rect 1468 1837 1470 1842
rect 1260 1827 1262 1831
rect 1282 1827 1284 1831
rect 1199 1806 1201 1811
rect 1374 1824 1376 1828
rect 1396 1824 1398 1828
rect 1261 1738 1263 1742
rect 1283 1738 1285 1742
rect 1400 1692 1402 1696
rect 1422 1692 1424 1696
rect 1779 1501 1781 1505
rect 1254 1495 1256 1499
rect 1276 1495 1278 1499
rect 880 1485 882 1489
rect 902 1485 904 1489
rect 1193 1474 1195 1479
rect 1368 1492 1370 1496
rect 1390 1492 1392 1496
rect 1801 1501 1803 1505
rect 1849 1502 1851 1506
rect 1045 1424 1047 1428
rect 1067 1424 1069 1428
rect 1093 1424 1096 1428
rect 1255 1406 1257 1410
rect 1277 1406 1279 1410
rect 885 1362 887 1366
rect 907 1362 909 1366
rect 1394 1360 1396 1364
rect 1416 1360 1418 1364
rect 825 1207 827 1212
rect 881 1206 883 1210
rect 903 1206 905 1210
rect 929 1206 932 1210
rect 1370 1158 1373 1167
<< ndiffusion >>
rect 1251 1802 1260 1803
rect 1256 1797 1260 1802
rect 1262 1799 1267 1803
rect 1272 1799 1282 1803
rect 1262 1797 1282 1799
rect 1284 1798 1298 1803
rect 1304 1798 1306 1803
rect 1466 1820 1468 1823
rect 1470 1820 1472 1823
rect 1476 1820 1478 1823
rect 1284 1797 1306 1798
rect 1365 1799 1374 1800
rect 1197 1789 1199 1792
rect 1201 1789 1203 1792
rect 1207 1789 1209 1792
rect 1370 1794 1374 1799
rect 1376 1796 1381 1800
rect 1386 1796 1396 1800
rect 1376 1794 1396 1796
rect 1398 1795 1412 1800
rect 1418 1795 1420 1800
rect 1398 1794 1420 1795
rect 1252 1710 1261 1711
rect 1257 1705 1261 1710
rect 1263 1707 1268 1711
rect 1273 1707 1283 1711
rect 1263 1705 1283 1707
rect 1285 1706 1299 1711
rect 1305 1706 1307 1711
rect 1285 1705 1307 1706
rect 1391 1667 1400 1668
rect 1396 1662 1400 1667
rect 1402 1664 1407 1668
rect 1412 1664 1422 1668
rect 1402 1662 1422 1664
rect 1424 1663 1438 1668
rect 1444 1663 1446 1668
rect 1424 1662 1446 1663
rect 1245 1470 1254 1471
rect 1250 1465 1254 1470
rect 1256 1467 1261 1471
rect 1266 1467 1276 1471
rect 1256 1465 1276 1467
rect 1278 1466 1292 1471
rect 1298 1466 1300 1471
rect 1770 1473 1779 1474
rect 1775 1468 1779 1473
rect 1781 1470 1786 1474
rect 1791 1470 1801 1474
rect 1781 1468 1801 1470
rect 1803 1469 1817 1474
rect 1823 1469 1824 1474
rect 1803 1468 1824 1469
rect 1836 1468 1839 1473
rect 1845 1468 1849 1473
rect 1851 1468 1854 1473
rect 1859 1468 1860 1473
rect 1278 1465 1300 1466
rect 1359 1467 1368 1468
rect 871 1457 880 1458
rect 876 1452 880 1457
rect 882 1454 887 1458
rect 892 1454 902 1458
rect 882 1452 902 1454
rect 904 1453 918 1458
rect 924 1453 926 1458
rect 1191 1457 1193 1460
rect 1195 1457 1197 1460
rect 1201 1457 1203 1460
rect 904 1452 926 1453
rect 1364 1462 1368 1467
rect 1370 1464 1375 1468
rect 1380 1464 1390 1468
rect 1370 1462 1390 1464
rect 1392 1463 1406 1468
rect 1412 1463 1414 1468
rect 1392 1462 1414 1463
rect 1036 1396 1045 1397
rect 1041 1391 1045 1396
rect 1047 1391 1067 1397
rect 1069 1391 1093 1397
rect 1096 1391 1101 1397
rect 1107 1391 1125 1397
rect 1246 1378 1255 1379
rect 1251 1373 1255 1378
rect 1257 1375 1262 1379
rect 1267 1375 1277 1379
rect 1257 1373 1277 1375
rect 1279 1374 1293 1379
rect 1299 1374 1301 1379
rect 1279 1373 1301 1374
rect 1385 1335 1394 1336
rect 876 1334 885 1335
rect 881 1329 885 1334
rect 887 1331 892 1335
rect 897 1331 907 1335
rect 887 1329 907 1331
rect 909 1330 923 1335
rect 929 1330 931 1335
rect 1390 1330 1394 1335
rect 1396 1332 1401 1336
rect 1406 1332 1416 1336
rect 1396 1330 1416 1332
rect 1418 1331 1432 1336
rect 1438 1331 1440 1336
rect 1418 1330 1440 1331
rect 909 1329 931 1330
rect 872 1178 881 1179
rect 820 1173 825 1178
rect 827 1173 831 1178
rect 838 1173 840 1178
rect 877 1173 881 1178
rect 883 1173 903 1179
rect 905 1173 929 1179
rect 932 1173 937 1179
rect 943 1173 961 1179
rect 1346 1109 1351 1118
rect 1361 1109 1370 1118
rect 1373 1109 1384 1118
rect 1395 1109 1399 1118
<< pdiffusion >>
rect 1460 1837 1461 1842
rect 1466 1837 1468 1842
rect 1470 1837 1472 1842
rect 1476 1837 1484 1842
rect 1258 1827 1260 1831
rect 1262 1827 1267 1831
rect 1272 1827 1282 1831
rect 1284 1827 1288 1831
rect 1293 1827 1294 1831
rect 1191 1806 1192 1811
rect 1197 1806 1199 1811
rect 1201 1806 1203 1811
rect 1207 1806 1215 1811
rect 1372 1824 1374 1828
rect 1376 1824 1381 1828
rect 1386 1824 1396 1828
rect 1398 1824 1402 1828
rect 1407 1824 1413 1828
rect 1259 1738 1261 1742
rect 1263 1738 1268 1742
rect 1273 1738 1283 1742
rect 1285 1738 1289 1742
rect 1398 1692 1400 1696
rect 1402 1692 1407 1696
rect 1412 1692 1422 1696
rect 1424 1692 1428 1696
rect 1433 1692 1439 1696
rect 1777 1501 1779 1505
rect 1781 1501 1786 1505
rect 1252 1495 1254 1499
rect 1256 1495 1261 1499
rect 1266 1495 1276 1499
rect 1278 1495 1282 1499
rect 1287 1495 1288 1499
rect 878 1485 880 1489
rect 882 1485 887 1489
rect 892 1485 902 1489
rect 904 1485 908 1489
rect 1185 1474 1186 1479
rect 1191 1474 1193 1479
rect 1195 1474 1197 1479
rect 1201 1474 1209 1479
rect 1366 1492 1368 1496
rect 1370 1492 1375 1496
rect 1380 1492 1390 1496
rect 1392 1492 1396 1496
rect 1401 1492 1407 1496
rect 1791 1501 1801 1505
rect 1803 1501 1807 1505
rect 1837 1502 1839 1506
rect 1844 1502 1849 1506
rect 1851 1502 1854 1506
rect 1859 1502 1860 1506
rect 1043 1424 1045 1428
rect 1047 1424 1052 1428
rect 1057 1424 1067 1428
rect 1069 1424 1073 1428
rect 1078 1424 1093 1428
rect 1096 1424 1101 1428
rect 1106 1424 1112 1428
rect 1253 1406 1255 1410
rect 1257 1406 1262 1410
rect 1267 1406 1277 1410
rect 1279 1406 1283 1410
rect 883 1362 885 1366
rect 887 1362 892 1366
rect 897 1362 907 1366
rect 909 1362 913 1366
rect 1392 1360 1394 1364
rect 1396 1360 1401 1364
rect 1406 1360 1416 1364
rect 1418 1360 1422 1364
rect 1427 1360 1433 1364
rect 813 1207 814 1212
rect 821 1207 825 1212
rect 827 1207 831 1212
rect 879 1206 881 1210
rect 883 1206 888 1210
rect 893 1206 903 1210
rect 905 1206 909 1210
rect 914 1206 929 1210
rect 932 1206 937 1210
rect 942 1206 948 1210
rect 1347 1158 1351 1167
rect 1361 1158 1370 1167
rect 1373 1158 1383 1167
rect 1394 1158 1399 1167
<< ndcontact >>
rect 1251 1797 1256 1802
rect 1267 1799 1272 1803
rect 1298 1798 1304 1803
rect 1462 1819 1466 1823
rect 1472 1819 1476 1823
rect 1193 1788 1197 1792
rect 1203 1788 1207 1792
rect 1365 1794 1370 1799
rect 1381 1796 1386 1800
rect 1412 1795 1418 1800
rect 1252 1705 1257 1710
rect 1268 1707 1273 1711
rect 1299 1706 1305 1711
rect 1391 1662 1396 1667
rect 1407 1664 1412 1668
rect 1438 1663 1444 1668
rect 1245 1465 1250 1470
rect 1261 1467 1266 1471
rect 1292 1466 1298 1471
rect 1770 1468 1775 1473
rect 1786 1470 1791 1474
rect 1817 1469 1823 1474
rect 1839 1468 1845 1473
rect 1854 1468 1859 1473
rect 871 1452 876 1457
rect 887 1454 892 1458
rect 918 1453 924 1458
rect 1187 1456 1191 1460
rect 1197 1456 1201 1460
rect 1359 1462 1364 1467
rect 1375 1464 1380 1468
rect 1406 1463 1412 1468
rect 1036 1391 1041 1396
rect 1101 1391 1107 1397
rect 1246 1373 1251 1378
rect 1262 1375 1267 1379
rect 1293 1374 1299 1379
rect 876 1329 881 1334
rect 892 1331 897 1335
rect 923 1330 929 1335
rect 1385 1330 1390 1335
rect 1401 1332 1406 1336
rect 1432 1331 1438 1336
rect 813 1173 820 1178
rect 831 1173 838 1178
rect 872 1173 877 1178
rect 937 1173 943 1179
rect 1351 1108 1361 1118
rect 1384 1109 1395 1119
<< pdcontact >>
rect 1461 1837 1466 1842
rect 1472 1837 1476 1842
rect 1253 1827 1258 1831
rect 1267 1827 1272 1831
rect 1288 1827 1293 1831
rect 1192 1806 1197 1811
rect 1203 1806 1207 1811
rect 1367 1824 1372 1828
rect 1381 1824 1386 1828
rect 1402 1824 1407 1828
rect 1254 1737 1259 1742
rect 1268 1737 1273 1742
rect 1289 1737 1294 1742
rect 1393 1692 1398 1696
rect 1407 1692 1412 1696
rect 1428 1692 1433 1696
rect 1772 1500 1777 1505
rect 1247 1495 1252 1499
rect 1261 1495 1266 1499
rect 1282 1495 1287 1499
rect 873 1484 878 1489
rect 887 1484 892 1489
rect 908 1484 913 1489
rect 1186 1474 1191 1479
rect 1197 1474 1201 1479
rect 1361 1492 1366 1496
rect 1375 1492 1380 1496
rect 1396 1492 1401 1496
rect 1786 1500 1791 1505
rect 1807 1500 1812 1505
rect 1839 1502 1844 1506
rect 1854 1502 1859 1506
rect 1038 1423 1043 1428
rect 1052 1423 1057 1428
rect 1073 1423 1078 1428
rect 1101 1423 1106 1428
rect 1248 1405 1253 1410
rect 1262 1405 1267 1410
rect 878 1361 883 1366
rect 892 1361 897 1366
rect 913 1361 918 1366
rect 1283 1405 1288 1410
rect 1387 1360 1392 1364
rect 1401 1360 1406 1364
rect 1422 1360 1427 1364
rect 814 1207 821 1212
rect 831 1207 838 1212
rect 874 1205 879 1210
rect 888 1205 893 1210
rect 909 1205 914 1210
rect 937 1205 942 1210
rect 1351 1158 1361 1168
rect 1383 1158 1394 1168
<< psubstratepcontact >>
rect 1263 1785 1269 1791
rect 1299 1785 1305 1791
rect 1377 1782 1383 1788
rect 1413 1782 1419 1788
rect 1264 1693 1270 1699
rect 1300 1693 1306 1699
rect 1403 1650 1409 1656
rect 1439 1650 1445 1656
rect 1257 1453 1263 1459
rect 1293 1453 1299 1459
rect 1371 1450 1377 1456
rect 1407 1450 1413 1456
rect 1782 1456 1788 1462
rect 1818 1456 1824 1462
rect 883 1440 889 1446
rect 919 1440 925 1446
rect 1048 1379 1054 1385
rect 1084 1379 1090 1385
rect 1258 1361 1264 1367
rect 1294 1361 1300 1367
rect 888 1317 894 1323
rect 924 1317 930 1323
rect 1397 1318 1403 1324
rect 1433 1318 1439 1324
rect 884 1161 890 1167
rect 920 1161 926 1167
<< nsubstratencontact >>
rect 1253 1838 1259 1843
rect 1288 1838 1293 1843
rect 1367 1835 1373 1840
rect 1402 1835 1407 1840
rect 1254 1746 1260 1751
rect 1289 1746 1294 1751
rect 1393 1703 1399 1708
rect 1428 1703 1433 1708
rect 873 1493 879 1498
rect 1247 1506 1253 1511
rect 1282 1506 1287 1511
rect 1772 1509 1778 1514
rect 1361 1503 1367 1508
rect 1396 1503 1401 1508
rect 1807 1509 1812 1514
rect 908 1493 913 1498
rect 1038 1432 1044 1437
rect 1073 1432 1078 1437
rect 878 1370 884 1375
rect 1248 1414 1254 1419
rect 1283 1414 1288 1419
rect 913 1370 918 1375
rect 1387 1371 1393 1376
rect 1422 1371 1427 1376
rect 874 1214 880 1219
rect 909 1214 914 1219
<< polysilicon >>
rect 1468 1842 1470 1845
rect 1260 1831 1262 1834
rect 1282 1831 1284 1834
rect 1374 1828 1376 1831
rect 1396 1828 1398 1831
rect 1468 1830 1470 1837
rect 1260 1819 1262 1827
rect 1199 1817 1262 1819
rect 1199 1811 1201 1817
rect 1199 1799 1201 1806
rect 1260 1803 1262 1817
rect 1282 1803 1284 1827
rect 1469 1826 1470 1830
rect 1374 1817 1376 1824
rect 1375 1811 1376 1817
rect 1200 1795 1201 1799
rect 1374 1800 1376 1811
rect 1396 1800 1398 1824
rect 1468 1823 1470 1826
rect 1468 1815 1470 1820
rect 1468 1810 1469 1815
rect 1199 1792 1201 1795
rect 1260 1793 1262 1797
rect 1199 1786 1201 1789
rect 1282 1777 1284 1797
rect 1374 1790 1376 1794
rect 1396 1792 1398 1794
rect 1396 1791 1452 1792
rect 1396 1790 1448 1791
rect 1282 1775 1285 1777
rect 1261 1742 1263 1745
rect 1283 1742 1285 1775
rect 1261 1728 1263 1738
rect 1262 1722 1263 1728
rect 1261 1711 1263 1722
rect 1283 1711 1285 1738
rect 1261 1701 1263 1705
rect 1283 1652 1285 1705
rect 1400 1696 1402 1699
rect 1422 1696 1424 1715
rect 1400 1685 1402 1692
rect 1401 1679 1402 1685
rect 1400 1668 1402 1679
rect 1422 1668 1424 1692
rect 1400 1658 1402 1662
rect 1422 1658 1424 1662
rect 1276 1649 1285 1652
rect 1276 1641 1278 1649
rect 1277 1636 1278 1641
rect 902 1536 903 1542
rect 880 1489 882 1492
rect 902 1489 904 1536
rect 1254 1499 1256 1502
rect 1276 1499 1278 1636
rect 1752 1528 1803 1531
rect 1779 1505 1781 1508
rect 1801 1505 1803 1528
rect 1849 1506 1851 1512
rect 1368 1496 1370 1499
rect 1390 1496 1392 1499
rect 880 1475 882 1485
rect 881 1469 882 1475
rect 880 1458 882 1469
rect 902 1458 904 1485
rect 1254 1487 1256 1495
rect 1193 1485 1256 1487
rect 1193 1479 1195 1485
rect 1193 1467 1195 1474
rect 1254 1471 1256 1485
rect 1276 1471 1278 1495
rect 1368 1485 1370 1492
rect 1369 1479 1370 1485
rect 1194 1463 1195 1467
rect 1368 1468 1370 1479
rect 1390 1468 1392 1492
rect 1779 1491 1781 1501
rect 1780 1485 1781 1491
rect 1779 1474 1781 1485
rect 1801 1474 1803 1501
rect 1849 1481 1851 1502
rect 1850 1477 1851 1481
rect 1849 1473 1851 1477
rect 1193 1460 1195 1463
rect 1254 1461 1256 1465
rect 1193 1454 1195 1457
rect 880 1400 882 1452
rect 902 1448 904 1452
rect 1276 1448 1278 1465
rect 1779 1464 1781 1468
rect 1801 1464 1803 1468
rect 1368 1458 1370 1462
rect 1390 1460 1392 1462
rect 1390 1459 1446 1460
rect 1390 1458 1442 1459
rect 1849 1461 1851 1468
rect 1276 1446 1279 1448
rect 1045 1428 1047 1431
rect 1067 1428 1069 1443
rect 1093 1428 1096 1442
rect 1045 1414 1047 1424
rect 908 1405 909 1412
rect 1046 1408 1047 1414
rect 795 1398 882 1400
rect 795 1220 797 1398
rect 885 1366 887 1369
rect 907 1366 909 1405
rect 1045 1397 1047 1408
rect 1067 1397 1069 1424
rect 1093 1397 1096 1424
rect 1255 1410 1257 1413
rect 1277 1410 1279 1446
rect 1255 1396 1257 1406
rect 1045 1387 1047 1391
rect 1067 1370 1069 1391
rect 1068 1366 1069 1370
rect 885 1352 887 1362
rect 886 1346 887 1352
rect 885 1335 887 1346
rect 907 1335 909 1362
rect 1093 1365 1096 1391
rect 1256 1390 1257 1396
rect 1255 1379 1257 1390
rect 1277 1379 1279 1406
rect 1255 1369 1257 1373
rect 1277 1369 1279 1373
rect 1095 1358 1096 1365
rect 1394 1364 1396 1367
rect 1416 1364 1418 1383
rect 1394 1353 1396 1360
rect 1395 1347 1396 1353
rect 1394 1336 1396 1347
rect 1416 1336 1418 1360
rect 885 1325 887 1329
rect 907 1325 909 1329
rect 1394 1326 1396 1330
rect 1416 1326 1418 1330
rect 795 1218 827 1220
rect 825 1212 827 1218
rect 881 1210 883 1213
rect 903 1210 905 1225
rect 929 1210 932 1224
rect 825 1178 827 1207
rect 881 1196 883 1206
rect 882 1190 883 1196
rect 881 1179 883 1190
rect 903 1179 905 1206
rect 929 1179 932 1206
rect 825 1169 827 1173
rect 881 1032 883 1173
rect 903 1133 905 1173
rect 929 1052 932 1173
rect 1370 1167 1373 1175
rect 1370 1140 1373 1158
rect 1370 1130 1371 1140
rect 1370 1118 1373 1130
rect 1370 1102 1373 1109
rect 929 1046 930 1052
rect 929 1038 932 1046
<< polycontact >>
rect 1465 1826 1469 1830
rect 1370 1811 1375 1817
rect 1196 1795 1200 1799
rect 1469 1810 1474 1815
rect 1448 1787 1452 1791
rect 1257 1722 1262 1728
rect 1422 1715 1426 1720
rect 1396 1679 1401 1685
rect 1272 1636 1277 1641
rect 903 1536 907 1542
rect 1743 1528 1752 1535
rect 876 1469 881 1475
rect 1364 1479 1369 1485
rect 1190 1463 1194 1467
rect 1775 1485 1780 1491
rect 1846 1477 1850 1481
rect 1442 1455 1446 1459
rect 904 1405 908 1412
rect 1041 1408 1046 1414
rect 1064 1366 1068 1370
rect 881 1346 886 1352
rect 1251 1390 1256 1396
rect 1416 1383 1420 1388
rect 1091 1358 1095 1365
rect 1390 1347 1395 1353
rect 877 1190 882 1196
rect 903 1127 908 1133
rect 1371 1130 1379 1140
rect 930 1046 938 1052
rect 881 1025 890 1032
<< metal1 >>
rect 768 1894 777 1897
rect 768 1890 1178 1894
rect 1498 1890 1508 1891
rect 768 1882 1508 1890
rect 768 1418 777 1882
rect 1096 1879 1508 1882
rect 1096 1878 1507 1879
rect 1440 1849 1458 1854
rect 925 1838 1253 1843
rect 1259 1838 1288 1843
rect 1293 1840 1305 1843
rect 1440 1840 1445 1849
rect 1462 1842 1466 1848
rect 1293 1838 1367 1840
rect 925 1837 1197 1838
rect 1193 1811 1197 1837
rect 845 1801 854 1802
rect 845 1799 1103 1801
rect 1203 1799 1207 1806
rect 845 1795 1196 1799
rect 845 1793 1103 1795
rect 1203 1794 1220 1799
rect 845 1594 854 1793
rect 1203 1792 1207 1794
rect 846 1475 853 1594
rect 882 1498 885 1764
rect 1193 1699 1197 1788
rect 1214 1728 1220 1794
rect 1231 1768 1235 1838
rect 1253 1831 1258 1838
rect 1288 1831 1293 1838
rect 1300 1835 1367 1838
rect 1373 1835 1402 1840
rect 1407 1835 1445 1840
rect 1367 1828 1372 1835
rect 1402 1828 1407 1835
rect 1472 1830 1476 1837
rect 1501 1831 1507 1878
rect 1487 1830 1507 1831
rect 1267 1816 1272 1827
rect 1267 1811 1318 1816
rect 1359 1811 1370 1817
rect 1267 1810 1363 1811
rect 1267 1805 1271 1810
rect 1267 1803 1272 1805
rect 1298 1803 1304 1810
rect 1315 1805 1363 1810
rect 1381 1807 1386 1824
rect 1402 1822 1407 1824
rect 1428 1826 1465 1830
rect 1428 1807 1432 1826
rect 1472 1825 1507 1830
rect 1472 1823 1476 1825
rect 1381 1802 1432 1807
rect 1381 1800 1386 1802
rect 1251 1791 1256 1797
rect 1412 1800 1418 1802
rect 1251 1785 1263 1791
rect 1269 1785 1299 1791
rect 1305 1785 1306 1791
rect 1365 1788 1370 1794
rect 1365 1782 1377 1788
rect 1383 1782 1413 1788
rect 1419 1782 1420 1788
rect 1231 1767 1275 1768
rect 1427 1767 1432 1802
rect 1231 1760 1410 1767
rect 1270 1751 1275 1760
rect 1260 1746 1289 1751
rect 1294 1746 1299 1751
rect 1256 1742 1259 1746
rect 1289 1742 1294 1746
rect 1214 1723 1257 1728
rect 1254 1722 1257 1723
rect 1268 1718 1273 1737
rect 1311 1718 1365 1719
rect 1268 1713 1365 1718
rect 1268 1711 1273 1713
rect 1299 1711 1305 1713
rect 1252 1699 1257 1705
rect 1193 1693 1264 1699
rect 1270 1693 1300 1699
rect 1306 1693 1307 1699
rect 1300 1655 1306 1693
rect 1358 1685 1365 1713
rect 1404 1708 1410 1760
rect 1422 1762 1432 1767
rect 1422 1720 1426 1762
rect 1399 1703 1428 1708
rect 1433 1703 1438 1708
rect 1393 1696 1398 1703
rect 1428 1696 1433 1703
rect 1358 1679 1396 1685
rect 1407 1675 1412 1692
rect 1428 1690 1433 1692
rect 1448 1675 1452 1787
rect 1407 1670 1452 1675
rect 1407 1668 1412 1670
rect 1438 1668 1444 1670
rect 1391 1656 1396 1662
rect 1391 1655 1403 1656
rect 1300 1650 1403 1655
rect 1409 1650 1439 1656
rect 1445 1655 1446 1656
rect 1462 1655 1466 1819
rect 1497 1815 1527 1818
rect 1474 1810 1527 1815
rect 1445 1650 1466 1655
rect 1321 1643 1328 1650
rect 1444 1649 1466 1650
rect 1258 1636 1272 1641
rect 1519 1564 1527 1810
rect 1519 1558 1752 1564
rect 907 1536 1495 1542
rect 1049 1506 1247 1511
rect 1253 1506 1282 1511
rect 1287 1508 1299 1511
rect 1287 1506 1361 1508
rect 1049 1502 1191 1506
rect 1049 1499 1055 1502
rect 919 1498 1055 1499
rect 879 1493 908 1498
rect 913 1493 1055 1498
rect 875 1489 878 1493
rect 908 1489 913 1493
rect 846 1470 876 1475
rect 846 1469 853 1470
rect 873 1469 876 1470
rect 887 1465 892 1484
rect 927 1465 950 1466
rect 998 1465 1006 1466
rect 887 1460 1006 1465
rect 887 1458 892 1460
rect 918 1458 924 1460
rect 927 1459 950 1460
rect 871 1446 876 1452
rect 978 1446 983 1447
rect 865 1440 883 1446
rect 889 1440 919 1446
rect 925 1440 983 1446
rect 767 1417 777 1418
rect 767 1412 776 1417
rect 767 1406 904 1412
rect 891 1375 897 1385
rect 978 1385 983 1440
rect 998 1415 1006 1460
rect 1049 1437 1055 1493
rect 1187 1479 1191 1502
rect 1154 1467 1163 1468
rect 1197 1467 1201 1474
rect 1154 1463 1190 1467
rect 1044 1432 1073 1437
rect 1078 1432 1083 1437
rect 1040 1428 1043 1432
rect 1073 1428 1078 1432
rect 998 1414 1036 1415
rect 998 1409 1041 1414
rect 1038 1408 1041 1409
rect 1052 1404 1057 1423
rect 1101 1404 1106 1423
rect 1052 1403 1106 1404
rect 1154 1403 1163 1463
rect 1197 1462 1214 1467
rect 1197 1460 1201 1462
rect 1052 1400 1163 1403
rect 1052 1399 1106 1400
rect 1101 1397 1106 1399
rect 1036 1385 1041 1391
rect 978 1379 1048 1385
rect 1054 1379 1084 1385
rect 1090 1381 1146 1385
rect 1090 1378 1147 1381
rect 884 1370 913 1375
rect 918 1370 923 1375
rect 880 1366 883 1370
rect 913 1366 918 1370
rect 1056 1366 1064 1370
rect 1136 1368 1147 1378
rect 1187 1368 1191 1456
rect 1208 1396 1214 1462
rect 1225 1436 1229 1506
rect 1247 1499 1252 1506
rect 1282 1499 1287 1506
rect 1294 1503 1361 1506
rect 1367 1503 1396 1508
rect 1401 1503 1406 1508
rect 1361 1496 1366 1503
rect 1396 1496 1401 1503
rect 1261 1484 1266 1495
rect 1261 1479 1312 1484
rect 1353 1479 1364 1485
rect 1261 1478 1357 1479
rect 1261 1473 1265 1478
rect 1261 1471 1266 1473
rect 1292 1471 1298 1478
rect 1309 1473 1357 1478
rect 1375 1475 1380 1492
rect 1396 1490 1401 1492
rect 1488 1476 1495 1536
rect 1423 1475 1495 1476
rect 1375 1470 1495 1475
rect 1375 1468 1380 1470
rect 1245 1459 1250 1465
rect 1406 1468 1412 1470
rect 1421 1469 1495 1470
rect 1245 1453 1257 1459
rect 1263 1453 1293 1459
rect 1299 1453 1300 1459
rect 1359 1456 1364 1462
rect 1359 1450 1371 1456
rect 1377 1450 1407 1456
rect 1413 1450 1414 1456
rect 1225 1435 1269 1436
rect 1421 1435 1426 1469
rect 1225 1428 1404 1435
rect 1264 1419 1269 1428
rect 1254 1414 1283 1419
rect 1288 1414 1293 1419
rect 1250 1410 1253 1414
rect 1283 1410 1288 1414
rect 1208 1391 1251 1396
rect 1248 1390 1251 1391
rect 1262 1386 1267 1405
rect 1305 1386 1359 1387
rect 1262 1381 1359 1386
rect 1262 1379 1267 1381
rect 1293 1379 1299 1381
rect 1136 1367 1192 1368
rect 1246 1367 1251 1373
rect 746 1353 757 1354
rect 745 1352 814 1353
rect 745 1345 881 1352
rect 746 1075 757 1345
rect 892 1342 897 1361
rect 1056 1342 1061 1366
rect 892 1337 1061 1342
rect 1079 1362 1085 1363
rect 1079 1358 1091 1362
rect 1136 1361 1258 1367
rect 1264 1361 1294 1367
rect 1300 1361 1301 1367
rect 892 1335 897 1337
rect 923 1335 929 1337
rect 876 1323 881 1329
rect 870 1317 888 1323
rect 894 1317 924 1323
rect 930 1317 1035 1323
rect 886 1219 892 1263
rect 854 1215 874 1219
rect 854 1212 858 1215
rect 880 1214 909 1219
rect 914 1214 919 1219
rect 838 1207 858 1212
rect 876 1210 879 1214
rect 909 1210 914 1214
rect 831 1196 838 1207
rect 831 1190 877 1196
rect 831 1178 838 1190
rect 888 1186 893 1205
rect 937 1186 942 1205
rect 1079 1186 1085 1358
rect 1139 1324 1149 1361
rect 1126 1317 1149 1324
rect 1294 1323 1300 1361
rect 1352 1353 1359 1381
rect 1398 1376 1404 1428
rect 1416 1430 1426 1435
rect 1416 1388 1420 1430
rect 1393 1371 1422 1376
rect 1427 1371 1432 1376
rect 1387 1364 1392 1371
rect 1422 1364 1427 1371
rect 1352 1347 1390 1353
rect 1401 1343 1406 1360
rect 1422 1358 1427 1360
rect 1442 1343 1446 1455
rect 1401 1338 1446 1343
rect 1463 1420 1472 1469
rect 1401 1336 1406 1338
rect 1432 1336 1438 1338
rect 1385 1324 1390 1330
rect 1385 1323 1397 1324
rect 1294 1318 1397 1323
rect 1403 1318 1433 1324
rect 1439 1318 1440 1324
rect 888 1182 1086 1186
rect 888 1181 942 1182
rect 1074 1181 1086 1182
rect 937 1179 942 1181
rect 813 1166 820 1173
rect 872 1167 877 1173
rect 866 1166 884 1167
rect 813 1161 884 1166
rect 890 1161 920 1167
rect 926 1166 927 1167
rect 1139 1166 1149 1317
rect 1349 1309 1358 1318
rect 1274 1182 1401 1194
rect 1463 1191 1473 1420
rect 1274 1181 1353 1182
rect 1383 1168 1393 1182
rect 926 1161 1150 1166
rect 813 1160 868 1161
rect 927 1159 1150 1161
rect 1351 1133 1360 1158
rect 1464 1140 1473 1191
rect 908 1127 1360 1133
rect 1379 1130 1473 1140
rect 1377 1129 1473 1130
rect 1455 1128 1473 1129
rect 1351 1118 1360 1127
rect 1329 1097 1371 1098
rect 1384 1097 1395 1109
rect 1329 1087 1398 1097
rect 1460 1075 1473 1128
rect 1519 1099 1527 1558
rect 1743 1535 1752 1558
rect 1787 1514 1795 1846
rect 1778 1509 1807 1514
rect 1812 1509 1844 1514
rect 1774 1505 1777 1509
rect 1807 1505 1812 1509
rect 1839 1506 1844 1509
rect 1583 1490 1775 1491
rect 1582 1486 1775 1490
rect 1582 1485 1766 1486
rect 1772 1485 1775 1486
rect 1582 1484 1763 1485
rect 746 1063 1473 1075
rect 746 1061 934 1063
rect 1467 1062 1473 1063
rect 1516 1053 1528 1099
rect 930 1052 1528 1053
rect 938 1046 1528 1052
rect 1516 1045 1528 1046
rect 1584 1034 1601 1484
rect 1786 1481 1791 1500
rect 1786 1477 1846 1481
rect 1786 1476 1824 1477
rect 1786 1474 1791 1476
rect 1817 1474 1823 1476
rect 1854 1473 1859 1502
rect 1770 1462 1775 1468
rect 1839 1462 1845 1468
rect 1764 1456 1782 1462
rect 1788 1456 1818 1462
rect 1824 1456 1845 1462
rect 1817 1276 1825 1456
rect 880 1032 1601 1034
rect 880 1025 881 1032
rect 890 1025 1601 1032
rect 1584 1023 1601 1025
<< m2contact >>
rect 916 1837 925 1843
rect 1458 1848 1466 1854
rect 882 1764 887 1769
rect 1787 1846 1796 1855
rect 1321 1633 1328 1643
rect 891 1385 897 1390
rect 1035 1317 1042 1323
rect 886 1263 892 1269
rect 1114 1317 1126 1324
rect 1349 1301 1358 1309
rect 1254 1180 1274 1197
rect 1319 1087 1329 1098
rect 1817 1261 1825 1276
<< metal2 >>
rect 1458 1854 1597 1855
rect 1466 1853 1597 1854
rect 1783 1853 1787 1854
rect 1466 1848 1787 1853
rect 1601 1846 1787 1848
rect 916 1772 924 1837
rect 916 1769 942 1772
rect 887 1764 942 1769
rect 934 1390 941 1764
rect 897 1385 941 1390
rect 935 1286 941 1385
rect 1321 1643 1328 1644
rect 1102 1323 1114 1324
rect 1042 1317 1114 1323
rect 1321 1312 1328 1633
rect 1319 1308 1329 1312
rect 1319 1302 1349 1308
rect 1257 1286 1273 1288
rect 935 1275 1273 1286
rect 935 1269 941 1275
rect 892 1263 942 1269
rect 1256 1197 1273 1275
rect 1319 1274 1329 1302
rect 1339 1301 1349 1302
rect 1319 1264 1817 1274
rect 1319 1098 1329 1264
rect 1825 1264 1826 1274
<< labels >>
rlabel metal1 1338 1652 1338 1652 1 Gnd
rlabel metal1 1313 1837 1313 1837 1 Vdd
rlabel metal1 848 1655 848 1655 1 in
rlabel metal1 1857 1488 1857 1488 7 out
rlabel metal1 1425 1805 1425 1805 1 Y
rlabel metal1 1426 1474 1426 1474 1 X
rlabel metal1 1264 1639 1264 1639 1 clk
<< end >>
