magic
tech scmos
timestamp 1608579289
<< nwell >>
rect 52 13 79 15
rect 221 13 248 15
rect -19 3 117 13
rect 150 3 286 13
rect 52 2 79 3
rect 221 2 248 3
<< polysilicon >>
rect 9 19 11 29
rect 178 19 180 29
rect -14 9 -12 11
rect -6 17 68 19
rect -6 9 -4 17
rect -2 9 0 11
rect 6 9 8 11
rect 14 9 16 11
rect 22 9 24 11
rect 26 9 28 17
rect 66 16 68 17
rect 33 9 35 11
rect 46 9 48 11
rect 58 9 60 11
rect 66 9 68 13
rect 74 9 76 11
rect 82 9 84 11
rect 104 9 106 11
rect -14 3 -12 6
rect -6 3 -4 6
rect -14 1 -4 3
rect -14 -19 -12 1
rect -6 -19 -4 1
rect -2 -19 0 6
rect 6 -5 8 6
rect 14 3 16 6
rect 22 3 24 6
rect 14 1 24 3
rect 6 -9 7 -5
rect 6 -19 8 -9
rect 14 -19 16 1
rect 22 -19 24 1
rect 26 -19 28 6
rect 33 -19 35 6
rect 46 -12 48 6
rect 58 -5 60 6
rect 46 -19 48 -16
rect 58 -19 60 -9
rect 66 -19 68 6
rect 155 9 157 11
rect 163 17 237 19
rect 163 9 165 17
rect 167 9 169 11
rect 175 9 177 11
rect 183 9 185 11
rect 191 9 193 11
rect 195 9 197 17
rect 235 16 237 17
rect 202 9 204 11
rect 215 9 217 11
rect 227 9 229 11
rect 235 9 237 13
rect 243 9 245 11
rect 251 9 253 11
rect 273 9 275 11
rect 74 -19 76 5
rect 82 2 84 5
rect 82 -19 84 -2
rect 104 -12 106 5
rect 104 -19 106 -16
rect 155 3 157 6
rect 163 3 165 6
rect 155 1 165 3
rect 155 -19 157 1
rect 163 -19 165 1
rect 167 -19 169 6
rect 175 -5 177 6
rect 183 3 185 6
rect 191 3 193 6
rect 183 1 193 3
rect 175 -9 176 -5
rect 175 -19 177 -9
rect 183 -19 185 1
rect 191 -19 193 1
rect 195 -19 197 6
rect 202 -19 204 6
rect 215 -12 217 6
rect 227 -5 229 6
rect 215 -19 217 -16
rect 227 -19 229 -9
rect 235 -19 237 6
rect 243 -19 245 5
rect 251 2 253 5
rect 251 -19 253 -2
rect 273 -12 275 5
rect 273 -19 275 -16
rect -14 -25 -12 -23
rect -6 -25 -4 -23
rect -2 -30 0 -23
rect 6 -25 8 -23
rect 14 -25 16 -23
rect 22 -30 24 -23
rect 26 -25 28 -23
rect 33 -25 35 -23
rect 46 -25 48 -23
rect 58 -25 60 -23
rect 66 -25 68 -23
rect 74 -30 76 -23
rect 82 -25 84 -23
rect 104 -25 106 -23
rect 155 -25 157 -23
rect -2 -32 76 -30
rect 163 -25 165 -23
rect 167 -30 169 -23
rect 175 -25 177 -23
rect 183 -25 185 -23
rect 191 -30 193 -23
rect 195 -25 197 -23
rect 202 -25 204 -23
rect 215 -25 217 -23
rect 227 -25 229 -23
rect 235 -25 237 -23
rect 243 -30 245 -23
rect 251 -25 253 -23
rect 273 -25 275 -23
rect 167 -32 245 -30
rect 27 -39 29 -32
rect 196 -39 198 -32
<< ndiffusion >>
rect 39 -19 44 -9
rect -15 -23 -14 -19
rect -12 -23 -11 -19
rect -7 -23 -6 -19
rect -4 -23 -2 -19
rect 0 -23 1 -19
rect 5 -23 6 -19
rect 8 -23 9 -19
rect 13 -23 14 -19
rect 16 -23 17 -19
rect 21 -23 22 -19
rect 24 -23 26 -19
rect 28 -23 33 -19
rect 35 -23 46 -19
rect 48 -23 58 -19
rect 60 -22 61 -19
rect 208 -19 213 -9
rect 65 -22 66 -19
rect 60 -23 66 -22
rect 68 -23 74 -19
rect 76 -23 77 -19
rect 81 -23 82 -19
rect 84 -23 87 -19
rect 91 -23 94 -19
rect 103 -23 104 -19
rect 106 -23 108 -19
rect 114 -23 116 -19
rect 154 -23 155 -19
rect 157 -23 158 -19
rect 162 -23 163 -19
rect 165 -23 167 -19
rect 169 -23 170 -19
rect 174 -23 175 -19
rect 177 -23 178 -19
rect 182 -23 183 -19
rect 185 -23 186 -19
rect 190 -23 191 -19
rect 193 -23 195 -19
rect 197 -23 202 -19
rect 204 -23 215 -19
rect 217 -23 227 -19
rect 229 -22 230 -19
rect 234 -22 235 -19
rect 229 -23 235 -22
rect 237 -23 243 -19
rect 245 -23 246 -19
rect 250 -23 251 -19
rect 253 -23 256 -19
rect 260 -23 263 -19
rect 272 -23 273 -19
rect 275 -23 277 -19
rect 283 -23 285 -19
rect -11 -32 -7 -23
rect 53 -26 57 -23
rect 69 -26 73 -23
rect 53 -29 73 -26
rect 158 -32 162 -23
rect 222 -26 226 -23
rect 238 -26 242 -23
rect 222 -29 242 -26
<< pdiffusion >>
rect -11 9 -7 19
rect -15 6 -14 9
rect -12 6 -6 9
rect -4 6 -2 9
rect 0 6 1 9
rect 5 6 6 9
rect 8 6 9 9
rect 13 6 14 9
rect 16 6 17 9
rect 53 13 66 16
rect 68 13 73 16
rect 53 9 57 13
rect 69 9 73 13
rect 21 6 22 9
rect 24 6 26 9
rect 28 6 33 9
rect 35 6 46 9
rect 48 6 58 9
rect 60 6 61 9
rect 65 6 66 9
rect 68 6 74 9
rect 69 5 74 6
rect 76 5 77 9
rect 81 5 82 9
rect 84 5 87 9
rect 91 5 94 9
rect 103 5 104 9
rect 106 5 108 9
rect 114 5 115 9
rect 158 9 162 19
rect 154 6 155 9
rect 157 6 163 9
rect 165 6 167 9
rect 169 6 170 9
rect 174 6 175 9
rect 177 6 178 9
rect 182 6 183 9
rect 185 6 186 9
rect 222 13 235 16
rect 237 13 242 16
rect 222 9 226 13
rect 238 9 242 13
rect 190 6 191 9
rect 193 6 195 9
rect 197 6 202 9
rect 204 6 215 9
rect 217 6 227 9
rect 229 6 230 9
rect 234 6 235 9
rect 237 6 243 9
rect 238 5 243 6
rect 245 5 246 9
rect 250 5 251 9
rect 253 5 256 9
rect 260 5 263 9
rect 272 5 273 9
rect 275 5 277 9
rect 283 5 284 9
<< metal1 >>
rect -19 24 61 26
rect 122 26 152 27
rect 65 24 230 26
rect 234 24 288 26
rect -19 19 -11 24
rect -7 20 17 24
rect 21 21 158 24
rect 21 20 103 21
rect -19 13 13 16
rect -19 10 -15 13
rect 9 10 13 13
rect 17 10 21 20
rect 29 11 38 15
rect 1 2 5 6
rect 1 -13 4 2
rect 29 -5 32 11
rect 61 9 65 20
rect 77 9 81 20
rect 98 9 103 20
rect 150 19 158 21
rect 162 20 186 24
rect 190 21 288 24
rect 190 20 272 21
rect 150 13 182 16
rect 150 10 154 13
rect 178 10 182 13
rect 186 10 190 20
rect 198 11 207 15
rect 11 -9 32 -5
rect 39 -2 80 1
rect 39 -5 44 -2
rect 53 -9 58 -5
rect 1 -16 46 -13
rect 50 -15 69 -12
rect 1 -19 5 -16
rect -19 -26 -15 -23
rect 9 -26 13 -23
rect -19 -29 13 -26
rect -19 -37 -11 -32
rect -7 -33 -3 -32
rect 17 -33 21 -23
rect 87 -19 91 5
rect 108 -2 114 5
rect 98 -16 102 -13
rect 109 -19 114 -6
rect 170 2 174 6
rect 170 -13 173 2
rect 198 -5 201 11
rect 230 9 234 20
rect 246 9 250 20
rect 267 9 272 20
rect 180 -9 201 -5
rect 208 -2 249 1
rect 208 -5 213 -2
rect 222 -9 227 -5
rect 170 -16 215 -13
rect 219 -15 238 -12
rect 170 -19 174 -16
rect 61 -33 65 -22
rect 77 -33 81 -23
rect 98 -33 103 -23
rect 150 -26 154 -23
rect 178 -26 182 -23
rect 150 -29 182 -26
rect -7 -37 3 -33
rect 7 -37 17 -33
rect 21 -37 61 -33
rect 65 -34 103 -33
rect 120 -34 158 -32
rect 65 -37 158 -34
rect 162 -33 166 -32
rect 186 -33 190 -23
rect 256 -19 260 5
rect 277 -2 283 5
rect 267 -16 271 -13
rect 278 -19 283 -2
rect 230 -33 234 -22
rect 246 -33 250 -23
rect 267 -33 272 -23
rect 162 -37 172 -33
rect 176 -37 186 -33
rect 190 -37 230 -33
rect 234 -34 272 -33
rect 234 -37 291 -34
rect 120 -38 152 -37
<< metal2 >>
rect 119 31 212 35
rect 38 24 43 30
rect 38 20 52 24
rect 38 16 43 20
rect 49 -5 52 20
rect 119 -2 122 31
rect 207 24 212 31
rect 207 20 221 24
rect 207 16 212 20
rect 39 -9 44 -5
rect 114 -6 122 -2
rect 218 -5 221 20
rect 208 -9 213 -5
rect 73 -16 94 -13
rect 98 -16 106 -13
rect 242 -16 263 -13
rect 267 -16 275 -13
<< ntransistor >>
rect -14 -23 -12 -19
rect -6 -23 -4 -19
rect -2 -23 0 -19
rect 6 -23 8 -19
rect 14 -23 16 -19
rect 22 -23 24 -19
rect 26 -23 28 -19
rect 33 -23 35 -19
rect 46 -23 48 -19
rect 58 -23 60 -19
rect 66 -23 68 -19
rect 74 -23 76 -19
rect 82 -23 84 -19
rect 104 -23 106 -19
rect 155 -23 157 -19
rect 163 -23 165 -19
rect 167 -23 169 -19
rect 175 -23 177 -19
rect 183 -23 185 -19
rect 191 -23 193 -19
rect 195 -23 197 -19
rect 202 -23 204 -19
rect 215 -23 217 -19
rect 227 -23 229 -19
rect 235 -23 237 -19
rect 243 -23 245 -19
rect 251 -23 253 -19
rect 273 -23 275 -19
<< ptransistor >>
rect -14 6 -12 9
rect -6 6 -4 9
rect -2 6 0 9
rect 6 6 8 9
rect 14 6 16 9
rect 66 13 68 16
rect 22 6 24 9
rect 26 6 28 9
rect 33 6 35 9
rect 46 6 48 9
rect 58 6 60 9
rect 66 6 68 9
rect 74 5 76 9
rect 82 5 84 9
rect 104 5 106 9
rect 155 6 157 9
rect 163 6 165 9
rect 167 6 169 9
rect 175 6 177 9
rect 183 6 185 9
rect 235 13 237 16
rect 191 6 193 9
rect 195 6 197 9
rect 202 6 204 9
rect 215 6 217 9
rect 227 6 229 9
rect 235 6 237 9
rect 243 5 245 9
rect 251 5 253 9
rect 273 5 275 9
<< polycontact >>
rect 7 -9 11 -5
rect 58 -9 62 -5
rect 46 -16 50 -12
rect 80 -2 84 2
rect 102 -16 106 -12
rect 176 -9 180 -5
rect 227 -9 231 -5
rect 215 -16 219 -12
rect 249 -2 253 2
rect 271 -16 275 -12
<< ndcontact >>
rect 39 -9 44 -5
rect -19 -23 -15 -19
rect -11 -23 -7 -19
rect 1 -23 5 -19
rect 9 -23 13 -19
rect 17 -23 21 -19
rect 61 -22 65 -18
rect 208 -9 213 -5
rect 77 -23 81 -19
rect 87 -23 91 -19
rect 98 -23 103 -19
rect 108 -23 114 -19
rect 150 -23 154 -19
rect 158 -23 162 -19
rect 170 -23 174 -19
rect 178 -23 182 -19
rect 186 -23 190 -19
rect 230 -22 234 -18
rect 246 -23 250 -19
rect 256 -23 260 -19
rect 267 -23 272 -19
rect 277 -23 283 -19
rect -11 -37 -7 -32
rect 158 -37 162 -32
<< pdcontact >>
rect -11 19 -7 24
rect 158 19 162 24
rect -19 6 -15 10
rect 1 6 5 10
rect 9 6 13 10
rect 17 6 21 10
rect 61 5 65 9
rect 77 5 81 9
rect 87 5 91 9
rect 98 5 103 9
rect 108 5 114 9
rect 150 6 154 10
rect 170 6 174 10
rect 178 6 182 10
rect 186 6 190 10
rect 230 5 234 9
rect 246 5 250 9
rect 256 5 260 9
rect 267 5 272 9
rect 277 5 283 9
<< m2contact >>
rect 38 11 43 16
rect 207 11 212 16
rect 49 -9 53 -5
rect 69 -16 73 -12
rect 109 -6 114 -2
rect 94 -16 98 -12
rect 218 -9 222 -5
rect 238 -16 242 -12
rect 263 -16 267 -12
<< psubstratepcontact >>
rect 61 24 65 28
rect 17 20 21 24
rect 230 24 234 28
rect 186 20 190 24
rect 3 -37 7 -33
rect 17 -37 21 -33
rect 61 -37 65 -33
rect 172 -37 176 -33
rect 186 -37 190 -33
rect 230 -37 234 -33
<< labels >>
rlabel polysilicon 28 -39 28 -39 1 b
rlabel polysilicon 10 28 10 28 5 a
rlabel metal1 -16 -35 -16 -35 2 Gnd
rlabel metal1 -16 21 -16 21 3 Vdd
rlabel metal1 90 -3 90 -3 1 f
rlabel polysilicon 179 28 179 28 1 a1
rlabel polysilicon 197 -39 197 -39 1 b1
rlabel metal1 259 -3 259 -3 1 f1
rlabel metal1 281 -4 281 -4 1 cout1
rlabel metal2 40 28 40 28 1 cin
<< end >>
