* SPICE3 file created from inv.ext - technology: scmos

M1000 f a Vdd w_n16_2# pmos w=5u l=2u
+  ad=30p pd=22u as=62p ps=54u
M1001 f a Gnd Gnd nmos w=4u l=2u
+  ad=28p pd=22u as=24p ps=20u
C0 w_n16_2# f 0.2fF
C1 a w_n16_2# 1.5fF
C2 Vdd w_n16_2# 0.8fF
C3 Gnd Gnd 1.9fF
C4 f Gnd 6.0fF
C5 a Gnd 9.8fF
C6 Vdd Gnd 2.1fF

VCC    Vdd     Gnd     DC=2.5


* The following two lines are for TRANSIENT analysis
*
*Vname +Node -Node Option T1  V1   T2  V2   T3   V3    T4  V4  T5   V5 
*----- ----- ----- ------ --  --   --  --   ---- --    --  --  ---- -- 
Vin     a     Gnd    PWL(   0   0    4N  0    4.1N 2.5   8N  2.5 8.1N  0  ) 


*     TSTEP TSTOP
*     ----- -----
.TRAN 0.1N  12N




* TEMPERATURE and OPTIONS SETTING

.OPTIONS TEMP=25 reltol = 1e-6 

*MODELS

.include tsmc_cmos025

.END
