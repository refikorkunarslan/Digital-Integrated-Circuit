* SPICE3 file created from nand2.ext - technology: scmos

M1000 f a Vdd Vdd pmos w=8u l=3u
+  ad=112p pd=44u as=80p ps=52u
M1001 Vdd b f Vdd pmos w=8u l=3u
+  ad=0p pd=0u as=0p ps=0u
M1002 a_14_13# a Gnd Gnd nmos w=8u l=3u
+  ad=80p pd=52u as=40p ps=26u
M1003 f b a_14_13# Gnd nmos w=8u l=3u
+  ad=40p pd=26u as=0p ps=0u
C0 Vdd a 4.9fF
C1 Vdd b 3.2fF
C2 Gnd a 3.2fF
C3 Vdd f 2.7fF
C4 Gnd b 8.6fF
C5 a b 0.3fF
C6 Gnd f 1.8fF
C7 Gnd a_14_13# 1.1fF
C8 b f 0.4fF

VCC    Vdd     Gnd     DC=2.5


* The following two lines are for TRANSIENT analysis
*
*Vname +Node -Node Option T1  V1   T2  V2   T3   V3    T4  V4  T5   V5 
*----- ----- ----- ------ --  --   --  --   ---- --    --  --  ---- -- 
Vin     a     Gnd    PWL(   0   0    4N  0    4.1N 2.5   8N  2.5 8.1N  0  ) 

* The following two lines are for TRANSIENT analysis
*
*Vname +Node -Node Option T1  V1   T2  V2   T3   V3    T4  V4  T5   V5 
*----- ----- ----- ------ --  --   --  --   ---- --    --  --  ---- -- 
Vi     b     Gnd    PWL(   0   0    4N  0    4.1N 2.5   8N  2.5 8.1N  0  ) 


*     TSTEP TSTOP
*     ----- -----
.TRAN 0.1N  12N


* The following line is for DC analysis

.DC VIN 0 2.6 0.1


* TEMPERATURE and OPTIONS SETTING

.OPTIONS TEMP=25 reltol = 1e-6 

*MODELS

.include tsmc_cmos025

.END
