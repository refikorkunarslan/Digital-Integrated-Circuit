* SPICE3 file created from nand2.ext - technology: scmos

.option scale=0.01u

M1000 f a Vdd Vdd pmos w=400 l=200
+  ad=800000 pd=4800 as=880000 ps=6000
M1001 Vdd b f Vdd pmos w=400 l=200
+  ad=0 pd=0 as=0 ps=0
M1002 f a Gnd Gnd nmos w=600 l=200
+  ad=2.52e+06 pd=10800 as=540000 ps=3000
M1003 f b f Gnd nmos w=600 l=200
+  ad=0 pd=0 as=0 ps=0
C0 Gnd Gnd 13.5fF
C1 f Gnd 14.2fF
C2 b Gnd 9.1fF
C3 a Gnd 9.1fF
C4 Vdd Gnd 2.1fF

VCC    Vdd     Gnd     DC=2.5


* The following two lines are for TRANSIENT analysis
*
*Vname +Node -Node Option T1  V1   T2  V2   T3   V3    T4  V4  T5   V5 
*----- ----- ----- ------ --  --   --  --   ---- --    --  --  ---- -- 
Vin     a     f    PWL(   0   0    4N  0    4.1N 2.5   8N  2.5 8.1N  0  ) 

* The following two lines are for TRANSIENT analysis
*
*Vname +Node -Node Option T1  V1   T2  V2   T3   V3    T4  V4  T5   V5 
*----- ----- ----- ------ --  --   --  --   ---- --    --  --  ---- -- 
Vi     b     f    PWL(   0   0    4N  0    4.1N 2.5   8N  2.5 8.1N  0  ) 

*     TSTEP TSTOP
*     ----- -----
.TRAN 0.1N  12N


* The following line is for DC analysis

.DC VIN 0 2.6 0.1


* TEMPERATURE and OPTIONS SETTING

.OPTIONS TEMP=25 reltol = 1e-6 

*MODELS

.include tsmc_cmos025

.END
