* SPICE3 file created from nor3.ext - technology: scmos

.option scale=1u

M1000 a_n4_4# a Vdd Vdd pmos w=4 l=2
+  ad=80 pd=48 as=28 ps=22
M1001 a_18_4# b a_n4_4# Vdd pmos w=4 l=2
+  ad=72 pd=44 as=0 ps=0
M1002 f c a_18_4# Vdd pmos w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1003 f a Gnd Gnd nmos w=6 l=2
+  ad=156 pd=76 as=162 ps=78
M1004 Gnd b f Gnd nmos w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1005 f c Gnd Gnd nmos w=6 l=2
+  ad=0 pd=0 as=0 ps=0
C0 Vdd f 0.4fF
C1 b f 0.2fF
C2 c Vdd 1.7fF
C3 a Vdd 1.7fF
C4 b Vdd 1.7fF
C5 c f 0.2fF
C6 Gnd Gnd 13.8fF
C7 f Gnd 11.8fF
C8 c Gnd 8.7fF
C9 b Gnd 9.1fF
C10 a Gnd 9.1fF

VCC    Vdd     Gnd     DC=2.5


* The following two lines are for TRANSIENT analysis
*
*Vname +Node -Node Option T1  V1   T2  V2   T3   V3    T4  V4  T5   V5 
*----- ----- ----- ------ --  --   --  --   ---- --    --  --  ---- -- 
Vin     a     f    PWL(   0   0    4N  0    4.1N 2.5   8N  2.5 8.1N  0  ) 

* The following two lines are for TRANSIENT analysis
*
*Vname +Node -Node Option T1  V1   T2  V2   T3   V3    T4  V4  T5   V5 
*----- ----- ----- ------ --  --   --  --   ---- --    --  --  ---- -- 
Vi     b     f    PWL(   0   0    4N  0    4.1N 2.5   8N  2.5 8.1N  0  ) 

* The following two lines are for TRANSIENT analysis
*
*Vname +Node -Node Option T1  V1   T2  V2   T3   V3    T4  V4  T5   V5 
*----- ----- ----- ------ --  --   --  --   ---- --    --  --  ---- -- 
V     c     f    PWL(   0   0    4N  0    4.1N 2.5   8N  2.5 8.1N  0  ) 

*     TSTEP TSTOP
*     ----- -----
.TRAN 0.1N  12N


* The following line is for DC analysis

.DC VIN 0 2.6 0.1


* TEMPERATURE and OPTIONS SETTING

.OPTIONS TEMP=25 reltol = 1e-6 

*MODELS

.include tsmc_cmos025

.END
